library verilog;
use verilog.vl_types.all;
entity Top_Level_vlg_vec_tst is
end Top_Level_vlg_vec_tst;
