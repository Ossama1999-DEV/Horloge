library verilog;
use verilog.vl_types.all;
entity cpt_dcpt_vlg_vec_tst is
end cpt_dcpt_vlg_vec_tst;
