library verilog;
use verilog.vl_types.all;
entity Afficheur_7_seg_vlg_vec_tst is
end Afficheur_7_seg_vlg_vec_tst;
